magic
tech scmos
timestamp 1637222525
<< error_p >>
rect 8 0 16 2
<< nwell >>
rect 5 5 30 28
<< ntransistor >>
rect 16 -5 18 -1
<< ptransistor >>
rect 16 14 18 22
<< ndiffusion >>
rect 15 -5 16 -1
rect 18 -5 19 -1
<< pdiffusion >>
rect 15 14 16 22
rect 18 14 19 22
<< ndcontact >>
rect 11 -5 15 -1
rect 19 -5 23 -1
<< pdcontact >>
rect 11 14 15 22
rect 19 14 23 22
<< polysilicon >>
rect 16 22 18 25
rect 16 -1 18 14
rect 16 -8 18 -5
<< polycontact >>
rect 12 0 16 4
<< metal1 >>
rect 5 27 30 31
rect 11 22 15 27
rect 19 4 23 14
rect 1 0 12 4
rect 19 0 39 4
rect 19 -1 23 0
rect 11 -9 15 -5
rect 4 -13 30 -9
<< labels >>
rlabel nwell 11 14 23 22 1 pdiff
rlabel nwell 5 5 30 8 1 VDD
rlabel space 11 -5 23 -1 1 ndiff
rlabel metal1 5 27 30 31 5 VDD
rlabel metal1 4 -13 30 -9 1 GND
rlabel metal1 1 0 16 4 1 INPUT
rlabel metal1 23 0 39 4 1 OUTPUT
<< end >>
